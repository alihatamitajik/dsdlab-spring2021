module uart (
    tx, rx, resetN, clk
);
    
endmodule