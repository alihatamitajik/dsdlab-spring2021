`timescale 1ns / 1ps

module tcam_tb;

endmodule