module processor (
    output [7:0] read_data,
    input [7:0] address,
    input write,
    input [7:0] write_data,
    input clk,
    input resetN
);
    
endmodule