module receiver(rx, rx_clk, [7:0] data_out, resetN, error, busy);
    
endmodule