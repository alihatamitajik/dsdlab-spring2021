module receiver(
    rx, 
    rx_clk, 
    [7:0] data_out, 
    resetN, 
    error, 
    busy);
    
    input rx, rx_clk, resetN;
    output data_out, error, busy;

    
endmodule 