module transmiter (tx, tx_clk, [7:0] data_in, start, busy, resetN);
    
endmodule