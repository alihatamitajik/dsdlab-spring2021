
module transmiter (tx, clk, tx_en, [7:0] data_in, start, busy, resetN);
    output reg tx, busy;
    input wire start, resetN, clk, rx_en, ;
    input [6:0] data_in;

    reg [7:0] data_send;
    reg [1:0] current_state = 0;
    reg [2:0] pos = 0;
    reg isStarted = 0;

    always @ (posedge clk or negedge resetN or posedge start) begin
        if (~resetN) begin                         // if module was reseted
            current_state <= 2b'00;                // go to Relax State
            isStarted <= 1b'0;                     // make not started
            tx <= 1b'1;                            // make tx 1
        end else if (start && ~isStarted) begin
            isStarted <= 1;                        // set started flag
            current_state <= 2b'01;                // Current State to Send Start Bit
            data_send <= {~^data_in,data_in};      // set data to send
        end else if (current_state == 2b'01) begin // If in Send Start Bit State
            if (tx_en) begin                       // If we are on rate
                tx <= 1b'0;                        // send start bit
                current_state <= 2b'10;            // go to next state - send data
            end
        end else if (current_state == 2b'10) begin // if in send data state
            if (tx_en) begin                       // if we are on rate
                tx <= data_send[pos];              // make tx the data in send position
                pos <= pos + 1;                    // add to position
                if (pos == 3b'111)begin            // if we reach position 7
                    current_state <= 2b'11         // go to next state - send stop bit
                end                  
            end 
        end else if (current_state == 2b'11) begin // if in send stop bit state
            if (tx_en) begin                       // if we are on rate
                tx <= 1b'1;                        // send stop bit (1)
                current_state <= 2b'00;            // go to relax state
            end
        end
    end
endmodule