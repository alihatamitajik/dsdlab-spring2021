module transmiter (
    tx, 
    tx_clk, 
    [6:0] data_in, 
    start, 
    busy, 
    resetN);

endmodule